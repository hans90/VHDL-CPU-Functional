entity SYSTEM is
end SYSTEM;

architecture FUNCTIONAL of SYSTEM is
begin


end architecture;

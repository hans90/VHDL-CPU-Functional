package body CPU_DEFS_PACK_BODY of CPU_DEFS_PACK is
begin
end CPU_DEFS_PACK_BODY;

package CPU_DEFS_PACK is
begin
end CPU_DEFS_PACK;
